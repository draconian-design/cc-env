{% include 'copyright' %}
{% set NAME = 'types' %}

`ifndef __{{ cookiecutter.package | upper }}_{{ NAME | upper }}_SV__
 `define __{{ cookiecutter.package | upper }}_{{ NAME | upper }}_SV__

`endif // guard
